module Element(input logic clk, reset,
												output logic y);

endmodule